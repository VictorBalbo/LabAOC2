library verilog;
use verilog.vl_types.all;
entity cache is
end cache;
