library verilog;
use verilog.vl_types.all;
entity RAM is
end RAM;
